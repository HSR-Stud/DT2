Y <= transport A or B after 9 ns;