variable var_name {, var_name}: type_name 
								[:= value];
