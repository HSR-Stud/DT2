Y <= inertial A or B after 9 ns;
--Achtung ist das gleiche:
Y <= A or B after 9 ns;