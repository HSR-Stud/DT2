entity <ENTITY_NAME> is
	port(
		{<PORT_NAME>: <mode> <type>;}
		);
end <ENTITY_NAME>;