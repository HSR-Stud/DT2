constant sym_cyc: time := 100 ns;