library <library_name> {,<libary_name>};
use <library_name>.<element_name>;	
--oder
use <library_name>.all			
--Beispiel
library ieee;
use ieee.std_logic_1164.all;