--Verwendung von Typenkonvertierung
Y <= To_StdLogicVector(A);
B <= To_bitvector(X);
