architecture <ARCHITECTURE_NAME> of <ENTITY_NAME> is
	-- Signaldeklerationen
	signal ....
	-- Komponentdeklerationen
	component ...
begin
	-- Anweisungsteil
end <ARCHITECTURE_NAME>;