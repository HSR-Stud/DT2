signal <sig_name> {, <sig_name>}: type;

Bsp: signal sig1, sig2: bit;
