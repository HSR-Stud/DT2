entity DEVICE is
	port(
		A, B: in bit_vector (3 downto 0);
		Y: out bit);
end DEVICE;