generic(param_name: param_type:=initial_value[;param_name: param_type:=initial_value]);