--Erfassen einer positiven Flanke 
--    des Signals CLK
if CLK'event and CLK = '1' then ...

--Erfassen einer negativen Flanke 
--    des Signals CLK
if CLK'event and CLK = '0' then ...
